library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DECO_INST is
    Port ( OPCODE : in  STD_LOGIC_VECTOR (4 downto 0);
           TIPOR : out  STD_LOGIC;
           BEQ : out  STD_LOGIC;
           BNEQ : out  STD_LOGIC;
           BLT : out  STD_LOGIC;
           BLE : out  STD_LOGIC;
           BGT : out  STD_LOGIC;
           BGET : out  STD_LOGIC
			 );
end DECO_INST;

architecture Behavioral of DECO_INST is
CONSTANT OPCODE_TIPOR 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
CONSTANT OPCODE_BEQI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01101";
CONSTANT OPCODE_BNEI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01110";
CONSTANT OPCODE_BLTI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01111";
CONSTANT OPCODE_BLETI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10000";
CONSTANT OPCODE_BGTI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10001";
CONSTANT OPCODE_BGETI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10010";
CONSTANT OPCODE_B			: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10011";

begin
	TIPOR <= '1' WHEN (OPCODE = OPCODE_TIPOR) ELSE '0';
	BEQ 	<= '1' WHEN (OPCODE = OPCODE_BEQI) ELSE '0';
	BNEQ 	<= '1' WHEN (OPCODE = OPCODE_BNEI) ELSE '0';
	BLT 	<= '1' WHEN (OPCODE = OPCODE_BLTI) ELSE '0';
	BLE 	<= '1' WHEN (OPCODE = OPCODE_BLETI) ELSE '0';
	BGT 	<= '1' WHEN (OPCODE = OPCODE_BGTI) ELSE '0';
	BGET	<= '1' WHEN (OPCODE = OPCODE_BGETI) ELSE '0';
end Behavioral;